;arr;arr_cp;length;eq;uniques;i;searchIndices;curr;return@NUL Array to make unique values only is passed in as arr;
CLR i;
ADD 0 -1 i;
LEN arr length;
SUB length 1 length;
NUL == Start Loop ==;
CLR searchIndices;
ADD i 1 i;
SWI length i 20;
LOD std::dup.spice ^arr arr_cp;
GET i arr_cp curr;
PUT 0 arr_cp curr;
LOD std::arrays\index_of.spice ^arr_cp searchIndices;
PUT 0 searchIndices i;
LOD std::math\equal.spice searchIndices eq;
NUL if searchIndices != i, skip adding;
SWI eq 1 6;
ADD 0 curr uniques;
SWI 0 1 6;
NUL == End Loop ==;
LOD std::dup.spice ^uniques return;