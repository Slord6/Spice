;target;result;@
ADD 0 0 target;
LOD fib.spice target result;
OUT result