;arr;val;tmp;maxI;i;compare;return@NUL arr set by caller. 0th element is value to find. Index returned offsets as if value to find wasn't present;
ADD 0 -1 return;
GET 0 arr val;
LEN arr tmp;
SUB tmp 1 maxI;
NUL;
NUL == Start Loop ==;
ADD 1 i i;
CLR compare;
CLR return;
CLR tmp;
ADD 0 val compare;
GET i arr compare;
LOD std::math\equal.spice compare tmp;
SUB i 1 return;
BRK 0 tmp tmp;
NUL if i < maxI goto line(8);
SWI i maxI 7;
NUL == END LOOP ==;
NUL Value not in array, return -1;
CLR return;
ADD 0 -1 return;