;x;return@
POW x 0.5 return;