;return@