;target;fib;fibEnd;r1;r2;count;fibLen;return;@
ALS // NUL;
// target is set to required # from LOD;
// Start we do manually;
ADD 0 0 fibLen;
PUT fibLen fib 0;
ADD 1 fibLen fibLen;
PUT fibLen fib 1;
ADD 1 fibLen fibLen;
PUT fibLen fib 1;
// LOOP START;
// Get last element in fib, store in r1;
GET fibLen fib r1;
// GET last-1 element in fib, store in r2;
SUB fibLen 1 r2;
GET r2 fib r2;
// Add elements, store in r1;
ADD r1 r2 r1;
// Increase tracked array index;
ADD 1 fibLen fibLen;
// Put new element in last position;
PUT fibLen fib r1;
OUT fib;
// Note - NUL (//) statements count towards line count, as does prog part 1, prior to '@';
SWI fibLen target 10;
// LOOP END;
// Get the target element and store in return;
GET target fib return;